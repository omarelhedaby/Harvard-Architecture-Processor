LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MEM_RTI_UNIT IS

	PORT (RTI_SIG, clk: IN STD_LOGIC;
    RTI_OUT: OUT STD_LOGIC
    );
END ENTITY MEM_RTI_UNIT;


ARCHITECTURE MEM_RTI_UNIT_ARCH OF MEM_RTI_UNIT IS
	SIGNAL Count : INTEGER RANGE 0 TO 7;

BEGIN	

	PROCESS(clk) IS
	BEGIN

		if FALLING_EDGE(clk) THEN
			IF (RTI_SIG = '1') AND (COUNT = 0) THEN
				Count <= Count + 1 ;
				RTI_OUT <= '1';
			ELSIF Count = 1 AND RTI_SIG = '0'  THEN
				Count <= 0;
				RTI_OUT <= '0';
			else
				RTI_OUT <= '0';	
			END IF;
		END IF;



	END PROCESS;     
END MEM_RTI_UNIT_ARCH;