LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY DU_REGISTER_FILE_CONTROL_UNIT IS 
	PORT ( WB_ENABLE : IN std_logic_vector (1 DOWNTO 0);
           WRITE_ADDRESS_1,WRITE_ADDRESS_2 : IN std_logic_vector (2 DOWNTO 0);
           WRITE_MUX_0,WRITE_MUX_1,WRITE_MUX_2,WRITE_MUX_3,WRITE_MUX_4,WRITE_MUX_5,WRITE_MUX_6,WRITE_MUX_7 : OUT std_logic;
           WRITE_EN_0,WRITE_EN_1,WRITE_EN_2,WRITE_EN_3,WRITE_EN_4,WRITE_EN_5,WRITE_EN_6,WRITE_EN_7 : OUT std_logic;
           WRITE_EN_0_IN,WRITE_EN_1_IN,WRITE_EN_2_IN,WRITE_EN_3_IN,WRITE_EN_4_IN,WRITE_EN_5_IN,WRITE_EN_6_IN,WRITE_EN_7_IN : IN std_logic
           );
END DU_REGISTER_FILE_CONTROL_UNIT;


ARCHITECTURE DU_REGISTER_FILE_CONTROL_UNIT_ARCH OF DU_REGISTER_FILE_CONTROL_UNIT is
    
    SIGNAL OR_ENABLES : STD_LOGIC;
    BEGIN
    
---------------------------------WRITE ENABLES PART
    OR_ENABLES <= '1' WHEN  (WRITE_EN_0_IN = '1' OR WRITE_EN_1_IN = '1' OR WRITE_EN_2_IN = '1' OR WRITE_EN_3_IN = '1' OR WRITE_EN_4_IN = '1' OR WRITE_EN_5_IN = '1' OR WRITE_EN_6_IN = '1' OR WRITE_EN_7_IN = '1') 
    ELSE '0';

    WRITE_EN_0 <= '1' WHEN (WRITE_ADDRESS_1 = "000" OR WRITE_ADDRESS_2 = "000") AND (WB_ENABLE = "01") AND (OR_ENABLES = '0')
    ELSE '1' WHEN (WRITE_ADDRESS_1 = "000" OR WRITE_ADDRESS_2 = "000") AND (WB_ENABLE = "10") 
    ELSE '0';

    
    WRITE_EN_1 <= '1' WHEN (WRITE_ADDRESS_1 = "001" OR WRITE_ADDRESS_2 = "001") AND (WB_ENABLE = "01") AND (OR_ENABLES = '0')
    ELSE '1' WHEN (WRITE_ADDRESS_1 = "001" OR WRITE_ADDRESS_2 = "001") AND (WB_ENABLE = "10") 
    ELSE '0';
    
    WRITE_EN_2 <= '1' WHEN (WRITE_ADDRESS_1 = "010" OR WRITE_ADDRESS_2 = "010") AND (WB_ENABLE = "01") AND (OR_ENABLES = '0')
    ELSE '1' WHEN (WRITE_ADDRESS_1 = "010" OR WRITE_ADDRESS_2 = "010") AND (WB_ENABLE = "10") 
    ELSE '0';
    
    WRITE_EN_3 <= '1' WHEN (WRITE_ADDRESS_1 = "011" OR WRITE_ADDRESS_2 = "011") AND (WB_ENABLE = "01") AND (OR_ENABLES = '0')
    ELSE '1' WHEN (WRITE_ADDRESS_1 = "011" OR WRITE_ADDRESS_2 = "011") AND (WB_ENABLE = "10") 
    ELSE '0';
    
    WRITE_EN_4 <= '1' WHEN (WRITE_ADDRESS_1 = "100" OR WRITE_ADDRESS_2 = "100") AND (WB_ENABLE = "01") AND (OR_ENABLES = '0')
    ELSE '1' WHEN (WRITE_ADDRESS_1 = "100" OR WRITE_ADDRESS_2 = "100") AND (WB_ENABLE = "10") 
    ELSE '0';
    
    WRITE_EN_5 <= '1' WHEN (WRITE_ADDRESS_1 = "101" OR WRITE_ADDRESS_2 = "101") AND (WB_ENABLE = "01") AND (OR_ENABLES = '0')
    ELSE '1' WHEN (WRITE_ADDRESS_1 = "101" OR WRITE_ADDRESS_2 = "101") AND (WB_ENABLE = "10") 
    ELSE '0';

    WRITE_EN_6 <= '1' WHEN (WRITE_ADDRESS_1 = "110" OR WRITE_ADDRESS_2 = "110") AND (WB_ENABLE = "01") AND (OR_ENABLES = '0')
    ELSE '1' WHEN (WRITE_ADDRESS_1 = "110" OR WRITE_ADDRESS_2 = "110") AND (WB_ENABLE = "10") 
    ELSE '0';
    
    WRITE_EN_7 <= '1' WHEN (WRITE_ADDRESS_1 = "111" OR WRITE_ADDRESS_2 = "111") AND (WB_ENABLE = "01") AND (OR_ENABLES = '0')
    ELSE '1' WHEN (WRITE_ADDRESS_1 = "111" OR WRITE_ADDRESS_2 = "111") AND (WB_ENABLE = "10") 
    ELSE '0';
-------------------------------------------------------MUXSE PART
 
    WRITE_MUX_0 <= '0' WHEN WRITE_ADDRESS_1 = "000"   
    ELSE '1' WHEN WRITE_ADDRESS_2 = "000"  
    ELSE '0';

    WRITE_MUX_1 <= '0' WHEN WRITE_ADDRESS_1 = "001"   
    ELSE '1' WHEN WRITE_ADDRESS_2 = "001"  
    ELSE '0';

    WRITE_MUX_2 <= '0' WHEN WRITE_ADDRESS_1 = "010"   
    ELSE '1' WHEN WRITE_ADDRESS_2 = "010"  
    ELSE '0';

    WRITE_MUX_3 <= '0' WHEN WRITE_ADDRESS_1 = "011"   
    ELSE '1' WHEN WRITE_ADDRESS_2 = "011"  
    ELSE '0';

    WRITE_MUX_4 <= '0' WHEN WRITE_ADDRESS_1 = "100"   
    ELSE '1' WHEN WRITE_ADDRESS_2 = "100"  
    ELSE '0';

    WRITE_MUX_5 <= '0' WHEN WRITE_ADDRESS_1 = "101"   
    ELSE '1' WHEN WRITE_ADDRESS_2 = "101"  
    ELSE '0';


    WRITE_MUX_6 <= '0' WHEN WRITE_ADDRESS_1 = "110"   
    ELSE '1' WHEN WRITE_ADDRESS_2 = "110"  
    ELSE '0';

    WRITE_MUX_7 <= '0' WHEN WRITE_ADDRESS_1 = "111"   
    ELSE '1' WHEN WRITE_ADDRESS_2 = "111"  
    ELSE '0';

END DU_REGISTER_FILE_CONTROL_UNIT_ARCH;
