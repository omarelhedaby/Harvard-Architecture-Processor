LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY	DU_HDU IS
	PORT
	( 
		HAZARD_EN : OUT std_logic; 
		OP1,OP2,INST_0_2_ID_EX_OUT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		ID_EX_MEM_READ : IN STD_LOGIC 
	);
END DU_HDU;

ARCHITECTURE DU_HDU_ARCH OF DU_HDU IS
BEGIN

PROCESS(OP1,OP2,INST_0_2_ID_EX_OUT,ID_EX_MEM_READ)
	BEGIN


	IF ((ID_EX_MEM_READ = '1') AND ((OP1 = INST_0_2_ID_EX_OUT ) OR (OP2 = INST_0_2_ID_EX_OUT ))) THEN
		HAZARD_EN<='1';
	ELSE 
		HAZARD_EN<='0';
	END IF;


END PROCESS;

END DU_HDU_ARCH;